 * �;�9���������*8@D gVägled bollen förbi alla hinder för att passera genom ringarna och öppna dörren till nästa nivå. �Använd knapp 4 för att flytta bollen åt vänster, knapp 6 för att flytta bollen åt höger och knapp 2 för att studsa med bollen. Se upp för taggiga föremål. ~Använd sugen för att krympa bollen och pumpen för att blåsa upp den igen. Stora bollar flyter på vatten men inte de små. |Samla kristaller för att få extrapoäng och lagra din spelposition. Samla kristallbollar för att ge din boll längre liv. aHopp och hastighetsökningar ökar dina krafter tillfälligt medan gummigolv ger dig extra studs. Tillbaka 
Bra gjort! 	Fortsätt Avsluta Bounce Spelet är slut Högsta poäng Anvisningar Nivå %U Du har klarat nivå %U! 	Nytt spel Nytt rekord! Nästa OK Paus